// set the timescale
`timescale 1 ns / 100 ps
module wtm_tb(); // testbenches take no arguments
 	// set up inputs of NAND gate as registers so they can be manipulated at will
 	reg [4:0]in1;
 	reg [4:0]in2;
 	
 	// clocks are useful for testbenches because they allow you to check your
 	// circuit at regular intervals large enough for signals to propagate
 	reg clock;
 	
 	// set up output of NAND gate as wire
	wire [6:0] out;
	wire [6:0] btest;
 	
 	// prepare any other variables you want - nothing is off-limits in a TB
 	integer num_errors;
 	
 	// instantiate the RCA
 	wtm test_wtm(in1, in2, out,btest);
 	
 	// begin simulation
 	initial begin
       	$display($time, " simulation start");
       	
       	clock = 1'b0;
       	
       	       	
   @(negedge clock);
       	in1 = 5'd2;
       	in2 = 5'd14;
			
	@(negedge clock); // wait for the clock to go negative
       	in1 = 5'd5;
       	in2 = 5'd16;
						
	@(negedge clock); // wait for the clock to go negative
       	in1 = 5'd17;
       	in2 = 5'd3;
			
   @(negedge clock);
	      $stop;
	   
 	end
 	
 	always
       	#10 clock = ~clock; // toggle clock every 10 timescale units
 	
endmodule
//module square(left,right,up,down,x,y,clk);
//input left,right,up,down,clk;
//output x,y;
//reg x,y;
//initial begin 
// x = 10'd0;
// y = 10'd0; 
//always @(posedge clk) begin 
// if(left) begin 
//	x <= x-1; 
// end 
// if(right) begin
//	x<=x+1;
// end
// if(up) begin
//	y<=y-1;
// end
// if(down) bein
//	y<=y+1;
// end
//end
//endmodule

	module and_gate#(parameter DATA_WIDTH=32)(
    input [DATA_WIDTH-1:0] INPUT_A,
	 input [DATA_WIDTH-1:0] INPUT_B,
    output [DATA_WIDTH-1:0] OUT_AB
    );
    generate
        genvar index;
        for(index=0;index<DATA_WIDTH;index=index+1'b1)
            begin: identifier_and
					 and (OUT_AB[index], INPUT_A[index], INPUT_B[index]);
            end
    endgenerate
endmodule